-------------------------------------------------------------------------------
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: Readout Control Module
-------------------------------------------------------------------------------
-- This file is part of 'kek_bpm_rfsoc_dev'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'kek_bpm_rfsoc_dev', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiLitePkg.all;

library work;
use work.AppPkg.all;

entity ReadoutCtrl is
   generic (
      TPD_G : time := 1 ns);
   port (
      -- DSP Interface
      dspClk          : in  sl;
      dspRst          : in  sl;
      sigGenTrig      : out slv(1 downto 0);
      ncoConfig       : out slv(31 downto 0);
      -- DAC Interface (dacClk domain)
      dacClk          : in  sl;
      dacRst          : in  sl;
      dacDbgEn        : out sl;
      dacIDbg         : out Slv48Array(NUM_DAC_CH_C-1 downto 0);
      dacQDbg         : out Slv48Array(NUM_DAC_CH_C-1 downto 0);
      -- AXI-Lite Interface
      axilClk         : in  sl;
      axilRst         : in  sl;
      axilReadMaster  : in  AxiLiteReadMasterType;
      axilReadSlave   : out AxiLiteReadSlaveType;
      axilWriteMaster : in  AxiLiteWriteMasterType;
      axilWriteSlave  : out AxiLiteWriteSlaveType);
end ReadoutCtrl;

architecture rtl of ReadoutCtrl is

   type RegType is record
      sigGenTrig     : slv(1 downto 0);
      ncoConfig      : slv(31 downto 0);
      dacDbgEn       : sl;
      dacIDbg        : Slv48Array(NUM_DAC_CH_C-1 downto 0);
      dacQDbg        : Slv48Array(NUM_DAC_CH_C-1 downto 0);
      axilReadSlave  : AxiLiteReadSlaveType;
      axilWriteSlave : AxiLiteWriteSlaveType;
   end record RegType;
   constant REG_INIT_C : RegType := (
      sigGenTrig     => (others => '0'),
      ncoConfig      => (others => '0'),
      dacDbgEn       => '1',
      dacIDbg        => (others => (others => '0')),
      dacQDbg        => (others => (others => '0')),
      axilReadSlave  => AXI_LITE_READ_SLAVE_INIT_C,
      axilWriteSlave => AXI_LITE_WRITE_SLAVE_INIT_C);

   signal r   : RegType := REG_INIT_C;
   signal rin : RegType;

begin

   comb : process (axilReadMaster, axilRst, axilWriteMaster, r) is
      variable v      : RegType;
      variable axilEp : AxiLiteEndPointType;
   begin
      -- Latch the current value
      v := r;

      -- Reset strobes
      v.sigGenTrig := (others => '0');

      ----------------------------------------------------------------------
      --                AXI-Lite Register Logic
      ----------------------------------------------------------------------

      -- Determine the transaction type
      axiSlaveWaitTxn(axilEp, axilWriteMaster, axilReadMaster, v.axilWriteSlave, v.axilReadSlave);

      -- Map the read registers
      axiSlaveRegister (axilEp, x"00", 0, v.sigGenTrig(0));  -- Live Display
      axiSlaveRegister (axilEp, x"04", 0, v.sigGenTrig(1));  -- Fault Buffering
      axiSlaveRegister (axilEp, x"08", 0, v.ncoConfig);  -- 32-bits, address: [0x8:0xB]
      -- Reserved: address: [0xC:0xF]

      axiSlaveRegister (axilEp, x"10", 0, v.dacDbgEn);
      axiSlaveRegister (axilEp, x"20", 0, v.dacIDbg(0));
      axiSlaveRegister (axilEp, x"28", 0, v.dacQDbg(0));
      axiSlaveRegister (axilEp, x"30", 0, v.dacIDbg(1));
      axiSlaveRegister (axilEp, x"38", 0, v.dacQDbg(1));

      -- Closeout the transaction
      axiSlaveDefault(axilEp, v.axilWriteSlave, v.axilReadSlave, AXI_RESP_DECERR_C);

      ----------------------------------------------------------------------

      -- Outputs
      axilWriteSlave <= r.axilWriteSlave;
      axilReadSlave  <= r.axilReadSlave;

      -- Reset
      if (axilRst = '1') then
         v := REG_INIT_C;
      end if;

      -- Register the variable for next clock cycle
      rin <= v;

   end process comb;

   seq : process (axilClk) is
   begin
      if rising_edge(axilClk) then
         r <= rin after TPD_G;
      end if;
   end process seq;

   U_sigGenTrig : entity surf.SynchronizerOneShotVector
      generic map(
         TPD_G   => TPD_G,
         WIDTH_G => 2)
      port map(
         clk     => dspClk,
         dataIn  => r.sigGenTrig,
         dataOut => sigGenTrig);

   U_ncoConfig : entity surf.SynchronizerVector
      generic map(
         TPD_G   => TPD_G,
         WIDTH_G => 32)
      port map(
         clk     => dspClk,
         dataIn  => r.ncoConfig,
         dataOut => ncoConfig);

   GEN_VEC :
   for i in NUM_DAC_CH_C-1 downto 0 generate

      U_dacIDbg : entity surf.SynchronizerVector
         generic map(
            TPD_G   => TPD_G,
            WIDTH_G => 48)
         port map(
            clk     => dacClk,
            dataIn  => r.dacIDbg(i),
            dataOut => dacIDbg(i));

      U_dacQDbg : entity surf.SynchronizerVector
         generic map(
            TPD_G   => TPD_G,
            WIDTH_G => 48)
         port map(
            clk     => dacClk,
            dataIn  => r.dacQDbg(i),
            dataOut => dacQDbg(i));

   end generate GEN_VEC;

   U_dacDbgEn : entity surf.Synchronizer
      generic map(
         TPD_G => TPD_G)
      port map(
         clk     => dacClk,
         dataIn  => r.dacDbgEn,
         dataOut => dacDbgEn);

end rtl;
